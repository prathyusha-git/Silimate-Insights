module design_logic_combo_1_13(input logic a,b,c, output logic y);
  assign y = (a & b) | c;
endmodule

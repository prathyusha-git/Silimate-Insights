module design_logic_combo_3_8(input logic a,b,c, output logic y);
  assign y = (a ^ b) ^ c;
endmodule

module design_logic_combo_1_27(input logic a,b,c, output logic y);
  assign y = (a & b) | c;
endmodule
